module ramControl(input clk,
		  input [9:0] xAddress,
		  input [8:0] yAddress,
		  inout data,
		  input w);
   
